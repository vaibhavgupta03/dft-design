// Designing a dft filter for N=4 by taking the first four points of the DFT matrix

module dft4point ( input wire clk, input wire reset, input wire start, input wire signed [15:0] x0, x1, x2, x3,
                  output reg signed [15:0] Xr [0:3],output reg signed [15:0] Xi [0:3] , output reg done);

input k,n;

reg signed [15:0] x[0:3];
reg signed [15:0] cosVal[0:3];
reg signed [15:0] sinVal[0:3];
reg signed [31:0] tempR, tempI;

always @(*) begin
  cosVal[0] = 16'sd32767; sinVal[0] = 16'sd0;
  cosVal[1] = 16'sd0; sinVal[1] = 16'sd32767;
  cosVal[2] = -16'sd32767; sinVal[2] = 16'sd0;
  cosVal[3] = 16'sd0; sinVal[3] = -16'sd32767;
end

always @(posedge clk or posedge reset) begin
  if (reset) begin
    done <= 1'b0;
    k<=0;
    n<=0;
    tempR <= 32'sd0;
    tempI <= 32'sd0;
  end
  else if (start) begin
    x[0] <= x0;
    x[1] <= x1;
    x[2] <= x2;
    x[3] <= x3;

    tempR <= 32'sd0;
    tempI <= 32'sd0;
    for (k = 0; k < 4; k = k + 1) begin
      tempR = 32'sd0;
      tempI = 32'sd0;
      for (n = 0; n < 4; n = n + 1) begin
        tempR = tempR + (x[n] * cosVal[(k*n)%4]);
        tempI = tempI - (x[n] * sinVal[(k*n)%4]);
      end
      Xr[k] <= tempR >>> 15; // Scaling down to fit in 16 bits
      Xi[k] <= tempI >>> 15; // Scaling down to fit in 16 bits
    end
    done <= 1'b1;
  end
end
endmodule
// Designing a dft filter for N=4 by taking the first four points of the DFT matrix

module dft4point ( input wire clk, input wire reset, input wire start, input wire signed [15:0] x0, x1, x2, x3,
                  output reg signed [15:0] Xr [0:3],output reg signed [15:0] Xi [0:3] , output reg done);
            

endmodule